module MAE (
    
);






endmodule