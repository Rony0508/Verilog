module weight_update(










);
/*---------------------------------------------------------------------------------*/

parameter N = 8;

/*---------------------------------------------------------------------------------*/
input 





/*---------------------------------------------------------------------------------*/
//go to weight_pref
output reg [N-1:0]





/*---------------------------------------------------------------------------------*/
//wire



//



//





/*---------------------------------------------------------------------------------*/








/*---------------------------------------------------------------------------------*/







/*---------------------------------------------------------------------------------*/











endmodule