module MSE (
    
);






endmodule