module input_pref();

/*---------------------------------------------------------------------------------*/
parameter N = 8;

/*---------------------------------------------------------------------------------*/
input en,clk,reset_n,buf_select;

input [N-1:0]pe11_in011,pe12_in012,pe13_in013,pe14_in014,pe15_in015,pe16_in016,pe17_in017,pe18_in018
,pe21_in021,pe22_in022,pe23_in023,pe24_in024,pe25_in025,pe26_in026,pe27_in027,pe28_in028
,pe31_in031,pe32_in032,pe33_in033,pe34_in034,pe35_in035,pe36_in036,pe37_in037,pe38_in038
,pe41_in041,pe42_in042,pe43_in043,pe44_in044,pe45_in045,pe46_in046,pe47_in047,pe48_in048;
/*---------------------------------------------------------------------------------*/
output




/*---------------------------------------------------------------------------------*/

/*---------------------------------------------------------------------------------*/
//擷取成8 bit fixed point







/*---------------------------------------------------------------------------------*/







/*---------------------------------------------------------------------------------*/











endmodule