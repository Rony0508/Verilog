module weight_pref(










);
/*---------------------------------------------------------------------------------*/

parameter N = 8;

/*---------------------------------------------------------------------------------*/
input en,clk,reset_n,buf_select;





/*---------------------------------------------------------------------------------*/
//go to SA
output reg [N-1:0]





/*---------------------------------------------------------------------------------*/
//wire



//



//





/*---------------------------------------------------------------------------------*/








/*---------------------------------------------------------------------------------*/







/*---------------------------------------------------------------------------------*/











endmodule