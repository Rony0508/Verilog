module GC_IN(sw_in,i011,i012,i013,i014,i015,i016,i017,i018,i021,i022,i023,i024,i025,i026,i027,i028,i031,i032,i033,i034,i035,i036,i037,i038,i041,i042,i043,i044,i045,i046,i047,i048
,i111,i112,i113,i114,i115,i116,i117,i118,i121,i122,i123,i124,i125,i126,i127,i128,i131,i132,i133,i134,i135,i136,i137,i138,i141,i142,i143,i144,i145,i146,i147,i148
,w011,w012,w013,w014,w015,w016,w017,w018,w021,w022,w023,w024,w025,w026,w027,w028,w031,w032,w033,w034,w035,w036,w037,w038,w041,w042,w043,w044,w045,w046,w047,w048
,w111,w112,w113,w114,w115,w116,w117,w118,w121,w122,w123,w124,w125,w126,w127,w128,w131,w132,w133,w134,w135,w136,w137,w138,w141,w142,w143,w144,w145,w146,w147,w148
,w211,w212,w213,w214,w215,w216,w217,w218,w221,w222,w223,w224,w225,w226,w227,w228,w231,w232,w233,w234,w235,w236,w237,w238,w241,w242,w243,w244,w245,w246,w247,w248
,lunda,gama,beta,select_m0,select_m1,select_m2,select_m3,select0,select1);
parameter N=8;

input [2:0]sw_in;

//Select and reset,clk
output reg select_m0,select_m1,select_m2,select_m3,select0,select1;

//Port
output reg[N-1:0]
//input
i011,i012,i013,i014,i015,i016,i017,i018,i021,i022,i023,i024,i025,i026,i027,i028,i031,i032,i033,i034,i035,i036,i037,i038,i041,i042,i043,i044,i045,i046,i047,i048
,i111,i112,i113,i114,i115,i116,i117,i118,i121,i122,i123,i124,i125,i126,i127,i128,i131,i132,i133,i134,i135,i136,i137,i138,i141,i142,i143,i144,i145,i146,i147,i148
//weight
,w011,w012,w013,w014,w015,w016,w017,w018,w021,w022,w023,w024,w025,w026,w027,w028,w031,w032,w033,w034,w035,w036,w037,w038,w041,w042,w043,w044,w045,w046,w047,w048
,w111,w112,w113,w114,w115,w116,w117,w118,w121,w122,w123,w124,w125,w126,w127,w128,w131,w132,w133,w134,w135,w136,w137,w138,w141,w142,w143,w144,w145,w146,w147,w148
,w211,w212,w213,w214,w215,w216,w217,w218,w221,w222,w223,w224,w225,w226,w227,w228,w231,w232,w233,w234,w235,w236,w237,w238,w241,w242,w243,w244,w245,w246,w247,w248;
output reg [2*N-1:0]lunda,gama,beta;
//output



always@(sw_in)
begin 
    case(sw_in)
	3'b000:
begin
select_m0=0;select_m1=0;select_m2=0;select_m3=0;select0=1;select1=0;
i011=1;i012=1;i013=1;i014=1;i015=1;i016=1;i017=1;i018=1;i021=1;i022=1;i023=1;i024=1;i025=1;i026=1;i027=1;i028=1;i031=1;i032=1;i033=1;i034=1;i035=1;i036=1;
i037=1;i038=1;i041=1;i042=1;i043=1;i044=1;i045=1;i046=1;i047=1;i048=1;i111=2;i112=2;i113=2;i114=2;i115=2;i116=2;i117=2;i118=2;i121=2;i122=2;i123=2;i124=2;
i125=2;i126=2;i127=2;i128=2;i131=2;i132=2;i133=2;i134=2;i135=2;i136=2;i137=2;i138=2;i141=2;i142=2;i143=2;i144=2;i145=2;i146=2;i147=2;i148=2;w011=3;w012=3;
w013=3;w014=3;w015=3;w016=3;w017=3;w018=3;w021=3;w022=3;w023=3;w024=3;w025=3;w026=3;w027=3;w028=3;w031=3;w032=3;w033=3;w034=3;w035=3;w036=3;w037=3;w038=3;
w041=3;w042=3;w043=3;w044=3;w045=3;w046=3;w047=3;w048=3;w111=4;w112=4;w113=4;w114=4;w115=4;w116=4;w117=4;w118=4;w121=4;w122=4;w123=4;w124=4;w125=4;w126=4;
w127=4;w128=4;w131=4;w132=4;w133=4;w134=4;w135=4;w136=4;w137=4;w138=4;w141=4;w142=4;w143=4;w144=4;w145=4;w146=4;w147=4;w148=4;w211=5;w212=5;w213=5;w214=5;
w215=5;w216=5;w217=5;w218=5;w221=5;w222=5;w223=5;w224=5;w225=5;w226=5;w227=5;w228=5;w231=5;w232=5;w233=5;w234=5;w235=5;w236=5;w237=5;w238=5;w241=5;w242=5;
w243=5;w244=5;w245=5;w246=5;w247=5;w248=5;lunda=2;gama=3;beta=4;
end

	3'b001:
begin
select_m0=0;select_m1=0;select_m2=0;select_m3=0;select0=1;select1=0;
i011=2;i012=2;i013=2;i014=2;i015=2;i016=2;i017=2;i018=2;i021=2;i022=2;i023=2;i024=2;i025=2;i026=2;i027=2;i028=2;i031=2;i032=2;i033=2;i034=2;i035=2;i036=2;
i037=2;i038=2;i041=2;i042=2;i043=2;i044=2;i045=2;i046=2;i047=2;i048=2;i111=1;i112=1;i113=1;i114=1;i115=1;i116=1;i117=1;i118=1;i121=1;i122=1;i123=1;i124=1;
i125=1;i126=1;i127=1;i128=1;i131=1;i132=1;i133=1;i134=1;i135=1;i136=1;i137=1;i138=1;i141=1;i142=1;i143=1;i144=1;i145=1;i146=1;i147=1;i148=1;w011=4;w012=4;
w013=4;w014=4;w015=4;w016=4;w017=4;w018=4;w021=4;w022=4;w023=4;w024=4;w025=4;w026=4;w027=4;w028=4;w031=4;w032=4;w033=4;w034=4;w035=4;w036=4;w037=4;w038=4;
w041=4;w042=4;w043=4;w044=4;w045=4;w046=4;w047=4;w048=4;w111=3;w112=3;w113=3;w114=3;w115=3;w116=3;w117=3;w118=3;w121=3;w122=3;w123=3;w124=3;w125=3;w126=3;
w127=3;w128=3;w131=3;w132=3;w133=3;w134=3;w135=3;w136=3;w137=3;w138=3;w141=3;w142=3;w143=3;w144=3;w145=3;w146=3;w147=3;w148=3;w211=2;w212=2;w213=2;w214=2;
w215=2;w216=2;w217=2;w218=2;w221=2;w222=2;w223=2;w224=2;w225=2;w226=2;w227=2;w228=2;w231=2;w232=2;w233=2;w234=2;w235=2;w236=2;w237=2;w238=2;w241=2;w242=2;
w243=2;w244=2;w245=2;w246=2;w247=2;w248=2;lunda=2;gama=3;beta=4;
end

	3'b010:
begin
select_m0=0;select_m1=0;select_m2=0;select_m3=0;select0=1;select1=0;
i011=3;i012=3;i013=3;i014=3;i015=3;i016=3;i017=3;i018=3;i021=3;i022=3;i023=3;i024=3;i025=3;i026=3;i027=3;i028=3;i031=3;i032=3;i033=3;i034=3;i035=3;i036=3;
i037=3;i038=3;i041=3;i042=3;i043=3;i044=3;i045=3;i046=3;i047=3;i048=3;i111=4;i112=4;i113=4;i114=4;i115=4;i116=4;i117=4;i118=4;i121=4;i122=4;i123=4;i124=4;
i125=4;i126=4;i127=4;i128=4;i131=4;i132=4;i133=4;i134=4;i135=4;i136=4;i137=4;i138=4;i141=4;i142=4;i143=4;i144=4;i145=4;i146=4;i147=4;i148=4;w011=2;w012=2;
w013=2;w014=2;w015=2;w016=2;w017=2;w018=2;w021=2;w022=2;w023=2;w024=2;w025=2;w026=2;w027=2;w028=2;w031=2;w032=2;w033=2;w034=2;w035=2;w036=2;w037=2;w038=2;
w041=2;w042=2;w043=2;w044=2;w045=2;w046=2;w047=2;w048=2;w111=5;w112=5;w113=5;w114=5;w115=5;w116=5;w117=5;w118=5;w121=5;w122=5;w123=5;w124=5;w125=5;w126=5;
w127=5;w128=5;w131=5;w132=5;w133=5;w134=5;w135=5;w136=5;w137=5;w138=5;w141=5;w142=5;w143=5;w144=5;w145=5;w146=5;w147=5;w148=5;w211=1;w212=1;w213=1;w214=1;
w215=1;w216=1;w217=1;w218=1;w221=1;w222=1;w223=1;w224=1;w225=1;w226=1;w227=1;w228=1;w231=1;w232=1;w233=1;w234=1;w235=1;w236=1;w237=1;w238=1;w241=1;w242=1;
w243=1;w244=1;w245=1;w246=1;w247=1;w248=1;lunda=2;gama=3;beta=4;
end
	3'b011:
begin
select_m0=0;select_m1=0;select_m2=0;select_m3=0;select0=1;select1=0;
i011=4;i012=4;i013=4;i014=4;i015=4;i016=4;i017=4;i018=4;i021=4;i022=4;i023=4;i024=4;i025=4;i026=4;i027=4;i028=4;i031=4;i032=4;i033=4;i034=4;i035=4;i036=4;
i037=4;i038=4;i041=4;i042=4;i043=4;i044=4;i045=4;i046=4;i047=4;i048=4;i111=1;i112=1;i113=1;i114=1;i115=1;i116=1;i117=1;i118=1;i121=1;i122=1;i123=1;i124=1;
i125=1;i126=1;i127=1;i128=1;i131=1;i132=1;i133=1;i134=1;i135=1;i136=1;i137=1;i138=1;i141=1;i142=1;i143=1;i144=1;i145=1;i146=1;i147=1;i148=1;w011=5;w012=5;
w013=5;w014=5;w015=5;w016=5;w017=5;w018=5;w021=5;w022=5;w023=5;w024=5;w025=5;w026=5;w027=5;w028=5;w031=5;w032=5;w033=5;w034=5;w035=5;w036=5;w037=5;w038=5;
w041=5;w042=5;w043=5;w044=5;w045=5;w046=5;w047=5;w048=5;w111=2;w112=2;w113=2;w114=2;w115=2;w116=2;w117=2;w118=2;w121=2;w122=2;w123=2;w124=2;w125=2;w126=2;
w127=2;w128=2;w131=2;w132=2;w133=2;w134=2;w135=2;w136=2;w137=2;w138=2;w141=2;w142=2;w143=2;w144=2;w145=2;w146=2;w147=2;w148=2;w211=3;w212=3;w213=3;w214=3;
w215=3;w216=3;w217=3;w218=3;w221=3;w222=3;w223=3;w224=3;w225=3;w226=3;w227=3;w228=3;w231=3;w232=3;w233=3;w234=3;w235=3;w236=3;w237=3;w238=3;w241=3;w242=3;
w243=3;w244=3;w245=3;w246=3;w247=3;w248=3;lunda=2;gama=3;beta=4;
end
	3'b100:
begin
select_m0=0;select_m1=0;select_m2=0;select_m3=0;select0=1;select1=0;
i011=2;i012=2;i013=2;i014=2;i015=2;i016=2;i017=2;i018=2;i021=2;i022=2;i023=2;i024=2;i025=2;i026=2;i027=2;i028=2;i031=2;i032=2;i033=2;i034=2;i035=2;i036=2;
i037=2;i038=2;i041=2;i042=2;i043=2;i044=2;i045=2;i046=2;i047=2;i048=2;i111=5;i112=5;i113=5;i114=5;i115=5;i116=5;i117=5;i118=5;i121=5;i122=5;i123=5;i124=5;
i125=5;i126=5;i127=5;i128=5;i131=5;i132=5;i133=5;i134=5;i135=5;i136=5;i137=5;i138=5;i141=5;i142=5;i143=5;i144=5;i145=5;i146=5;i147=5;i148=5;w011=4;w012=4;
w013=4;w014=4;w015=4;w016=4;w017=4;w018=4;w021=4;w022=4;w023=4;w024=4;w025=4;w026=4;w027=4;w028=4;w031=4;w032=4;w033=4;w034=4;w035=4;w036=4;w037=4;w038=4;
w041=4;w042=4;w043=4;w044=4;w045=4;w046=4;w047=4;w048=4;w111=3;w112=3;w113=3;w114=3;w115=3;w116=3;w117=3;w118=3;w121=3;w122=3;w123=3;w124=3;w125=3;w126=3;
w127=3;w128=3;w131=3;w132=3;w133=3;w134=3;w135=3;w136=3;w137=3;w138=3;w141=3;w142=3;w143=3;w144=3;w145=3;w146=3;w147=3;w148=3;w211=1;w212=1;w213=1;w214=1;
w215=1;w216=1;w217=1;w218=1;w221=1;w222=1;w223=1;w224=1;w225=1;w226=1;w227=1;w228=1;w231=1;w232=1;w233=1;w234=1;w235=1;w236=1;w237=1;w238=1;w241=1;w242=1;
w243=1;w244=1;w245=1;w246=1;w247=1;w248=1;lunda=2;gama=3;beta=4;
end
	3'b101:
begin
select_m0=0;select_m1=0;select_m2=0;select_m3=0;select0=1;select1=0;
i011=3;i012=3;i013=3;i014=3;i015=3;i016=3;i017=3;i018=3;i021=3;i022=3;i023=3;i024=3;i025=3;i026=3;i027=3;i028=3;i031=3;i032=3;i033=3;i034=3;i035=3;i036=3;
i037=3;i038=3;i041=3;i042=3;i043=3;i044=3;i045=3;i046=3;i047=3;i048=3;i111=2;i112=2;i113=2;i114=2;i115=2;i116=2;i117=2;i118=2;i121=2;i122=2;i123=2;i124=2;
i125=2;i126=2;i127=2;i128=2;i131=2;i132=2;i133=2;i134=2;i135=2;i136=2;i137=2;i138=2;i141=2;i142=2;i143=2;i144=2;i145=2;i146=2;i147=2;i148=2;w011=1;w012=1;
w013=1;w014=1;w015=1;w016=1;w017=1;w018=1;w021=1;w022=1;w023=1;w024=1;w025=1;w026=1;w027=1;w028=1;w031=1;w032=1;w033=1;w034=1;w035=1;w036=1;w037=1;w038=1;
w041=1;w042=1;w043=1;w044=1;w045=1;w046=1;w047=1;w048=1;w111=5;w112=5;w113=5;w114=5;w115=5;w116=5;w117=5;w118=5;w121=5;w122=5;w123=5;w124=5;w125=5;w126=5;
w127=5;w128=5;w131=5;w132=5;w133=5;w134=5;w135=5;w136=5;w137=5;w138=5;w141=5;w142=5;w143=5;w144=5;w145=5;w146=5;w147=5;w148=5;w211=4;w212=4;w213=4;w214=4;
w215=4;w216=4;w217=4;w218=4;w221=4;w222=4;w223=4;w224=4;w225=4;w226=4;w227=4;w228=4;w231=4;w232=4;w233=4;w234=4;w235=4;w236=4;w237=4;w238=4;w241=4;w242=4;
w243=4;w244=4;w245=4;w246=4;w247=4;w248=4;lunda=2;gama=3;beta=4;
end
	3'b110:
begin
select_m0=0;select_m1=0;select_m2=0;select_m3=0;select0=1;select1=0;
i011=5;i012=5;i013=5;i014=5;i015=5;i016=5;i017=5;i018=5;i021=5;i022=5;i023=5;i024=5;i025=5;i026=5;i027=5;i028=5;i031=5;i032=5;i033=5;i034=5;i035=5;i036=5;
i037=5;i038=5;i041=5;i042=5;i043=5;i044=5;i045=5;i046=5;i047=5;i048=5;i111=1;i112=1;i113=1;i114=1;i115=1;i116=1;i117=1;i118=1;i121=1;i122=1;i123=1;i124=1;
i125=1;i126=1;i127=1;i128=1;i131=1;i132=1;i133=1;i134=1;i135=1;i136=1;i137=1;i138=1;i141=1;i142=1;i143=1;i144=1;i145=1;i146=1;i147=1;i148=1;w011=2;w012=2;
w013=2;w014=2;w015=2;w016=2;w017=2;w018=2;w021=2;w022=2;w023=2;w024=2;w025=2;w026=2;w027=2;w028=2;w031=2;w032=2;w033=2;w034=2;w035=2;w036=2;w037=2;w038=2;
w041=2;w042=2;w043=2;w044=2;w045=2;w046=2;w047=2;w048=2;w111=4;w112=4;w113=4;w114=4;w115=4;w116=4;w117=4;w118=4;w121=4;w122=4;w123=4;w124=4;w125=4;w126=4;
w127=4;w128=4;w131=4;w132=4;w133=4;w134=4;w135=4;w136=4;w137=4;w138=4;w141=4;w142=4;w143=4;w144=4;w145=4;w146=4;w147=4;w148=4;w211=3;w212=3;w213=3;w214=3;
w215=3;w216=3;w217=3;w218=3;w221=3;w222=3;w223=3;w224=3;w225=3;w226=3;w227=3;w228=3;w231=3;w232=3;w233=3;w234=3;w235=3;w236=3;w237=3;w238=3;w241=3;w242=3;
w243=3;w244=3;w245=3;w246=3;w247=3;w248=3;lunda=2;gama=3;beta=4;
end
	default:
begin
select_m0=0;select_m1=0;select_m2=0;select_m3=0;select0=1;select1=0;
i011=3;i012=3;i013=3;i014=3;i015=3;i016=3;i017=3;i018=3;i021=3;i022=3;i023=3;i024=3;i025=3;i026=3;i027=3;i028=3;i031=3;i032=3;i033=3;i034=3;i035=3;i036=3;
i037=3;i038=3;i041=3;i042=3;i043=3;i044=3;i045=3;i046=3;i047=3;i048=3;i111=5;i112=5;i113=5;i114=5;i115=5;i116=5;i117=5;i118=5;i121=5;i122=5;i123=5;i124=5;
i125=5;i126=5;i127=5;i128=5;i131=5;i132=5;i133=5;i134=5;i135=5;i136=5;i137=5;i138=5;i141=5;i142=5;i143=5;i144=5;i145=5;i146=5;i147=5;i148=5;w011=4;w012=4;
w013=4;w014=4;w015=4;w016=4;w017=4;w018=4;w021=4;w022=4;w023=4;w024=4;w025=4;w026=4;w027=4;w028=4;w031=4;w032=4;w033=4;w034=4;w035=4;w036=4;w037=4;w038=4;
w041=4;w042=4;w043=4;w044=4;w045=4;w046=4;w047=4;w048=4;w111=1;w112=1;w113=1;w114=1;w115=1;w116=1;w117=1;w118=1;w121=1;w122=1;w123=1;w124=1;w125=1;w126=1;
w127=1;w128=1;w131=1;w132=1;w133=1;w134=1;w135=1;w136=1;w137=1;w138=1;w141=1;w142=1;w143=1;w144=1;w145=1;w146=1;w147=1;w148=1;w211=2;w212=2;w213=2;w214=2;
w215=2;w216=2;w217=2;w218=2;w221=2;w222=2;w223=2;w224=2;w225=2;w226=2;w227=2;w228=2;w231=2;w232=2;w233=2;w234=2;w235=2;w236=2;w237=2;w238=2;w241=2;w242=2;
w243=2;w244=2;w245=2;w246=2;w247=2;w248=2;lunda=2;gama=3;beta=4;
end
    endcase
end

endmodule
